# BSD 3-Clause License
#
# Copyright 2024 Piyush Kumar, Da Eun Shim, Dongwon Jang, Azad Naeemi, or Georgia Institute of Technology
#
# Redistribution and use in source and binary forms, with or without 
# modification, are permitted provided that the following conditions are met:
#
# 1. Redistributions of source code must retain the above copyright notice, 
# this list of conditions and the following disclaimer.
#
# 2. Redistributions in binary form must reproduce the above copyright notice, 
# this list of conditions and the following disclaimer in the documentation 
# and/or other materials provided with the distribution.
#
# 3. Neither the name of the copyright holder nor the names of its contributors 
# may be used to endorse or promote products derived from this software without 
# specific prior written permission.
#
# THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS “AS IS” 
# AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, 
# THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE 
# ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE 
# FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES 
# (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; 
# LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND 
# ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT 
# (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS 
# SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.


VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.0005 ;

PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
  LAYER LEF58_PITCH STRING ;
  LAYER LEF58_GAP STRING ;
  LAYER LEF58_EOLKEEPOUT STRING ;
  LAYER LEF58_SPACING STRING ;
  LAYER LEF58_CORNERSPACING STRING ;
  LAYER LEF58_WIDTHTABLE STRING ;
  LAYER LEF58_CUTCLASS STRING ;
  LAYER LEF58_SPACINGTABLE STRING ;
  LAYER LEF58_ENCLOSURE STRING ;
  LAYER LEF58_RIGHTWAYONGRIDONLY STRING ;
  LAYER LEF58_RECTONLY STRING ;
END PROPERTYDEFINITIONS

LAYER BPR
  TYPE MASTERSLICE ;
END BPR

LAYER NW
  TYPE MASTERSLICE ;
END NW

LAYER ACT
  TYPE MASTERSLICE ;
END ACT

LAYER CONT
  TYPE MASTERSLICE ;
END CONT

LAYER GATE
  TYPE MASTERSLICE ;
END GATE

LAYER DUMMY
  TYPE MASTERSLICE ;
END DUMMY

LAYER NIM
  TYPE MASTERSLICE ;
END NIM

LAYER PIM
  TYPE MASTERSLICE ;
END PIM

LAYER SDCON
  TYPE MASTERSLICE ;
END SDCON

LAYER VBPR
  TYPE CUT ;
  SPACING 0.012 ;
  WIDTH 0.012 ;
END VBPR

LAYER VSD
  TYPE CUT ;
  SPACING 0.012 ;
  WIDTH 0.012 ;
END VSD

LAYER VG
  TYPE CUT ;
  SPACING 0.012 ;
  WIDTH 0.012 ;
END VG

LAYER M0
  TYPE ROUTING ;
  SPACING 0.012 ;
  WIDTH 0.012 ;
  PITCH 0.024 ;
  OFFSET 0.024 ;
  AREA 0.000288 ;
  MINSIZE 0.024 0.012 ;
  DIRECTION HORIZONTAL  ;
  PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.015 EXTENSION 0 0 0.017 ;" ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER CORNERTOCORNER WIDTH 0.000 SPACING 0.015 ; " ;
  PROPERTY LEF58_RECTONLY "RECTONLY ;" ;
END M0

LAYER V0
  TYPE CUT ;
  SPACING 0.012 ;
  WIDTH 0.012 ;
END V0

LAYER M1
  TYPE ROUTING ;
  SPACING 0.014 ;
  WIDTH 0.014 ;
  PITCH 0.042 ;
  OFFSET 0.021 ;
  AREA 0.000392 ;
  MINSIZE 0.014 0.028 ;
  DIRECTION VERTICAL ;
  PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.016 EXTENSION 0 0 0.020 ;" ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER CORNERTOCORNER WIDTH 0.000 SPACING 0.016 ; " ;
  PROPERTY LEF58_RECTONLY "RECTONLY ;" ;
END M1

LAYER V1
  TYPE CUT ;
  SPACING 0.012 ;
  WIDTH 0.012 ;
  ENCLOSURE BELOW 0.004 0 ;
  ENCLOSURE ABOVE 0.004 0 ;
END V1

LAYER M2
  TYPE ROUTING ;
  SPACING 0.012 ;
  SPACING 0.012 SAMENET ;
  WIDTH 0.012 ;
  PITCH 0.024 ;
  OFFSET 0.024 ;
  AREA 0.000288 ;
  MINSIZE 0.024 0.012 ;
  DIRECTION HORIZONTAL ;
  PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.015 EXTENSION 0 0 0.017 ;" ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER CORNERTOCORNER WIDTH 0.000 SPACING 0.015 ; " ;
  PROPERTY LEF58_RECTONLY "RECTONLY ;" ;
END M2

LAYER V2
  TYPE CUT ;
  SPACING 0.012 ;
  WIDTH 0.012 ;
  ENCLOSURE BELOW 0.004 0 ;
  ENCLOSURE ABOVE 0.004 0 ;
END V2

LAYER M3
  TYPE ROUTING ;
  SPACING 0.014 ;
  SPACING 0.014 SAMENET ;
  WIDTH 0.014 ;
  PITCH 0.028 ;
  AREA 0.000392 ;
  MINSIZE 0.014 0.028 ;
  DIRECTION VERTICAL ;
  PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.015 EXTENSION 0 0 0.020 ;" ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER CORNERTOCORNER WIDTH 0.000 SPACING 0.016 ; " ;
  PROPERTY LEF58_RECTONLY "RECTONLY ;" ;
END M3

LAYER V3
  TYPE CUT ;
  SPACING 0.014 ;
  WIDTH 0.014 ;
  ENCLOSURE BELOW 0.004 0 ;
  ENCLOSURE ABOVE 0.004 0 ;
END V3

LAYER M4
  TYPE ROUTING ;
  SPACING 0.021 ;
  SPACING 0.021 SAMENET ;
  WIDTH 0.021 ;
  PITCH 0.042 ;
  AREA 0.000882 ;
  MINSIZE 0.042 0.021 ;
  DIRECTION HORIZONTAL ;
  PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.022 EXTENSION 0 0 0.030 ;" ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER CORNERTOCORNER WIDTH 0.000 SPACING 0.024 ; " ;
  PROPERTY LEF58_RECTONLY "RECTONLY ;" ;
END M4

LAYER V4
  TYPE CUT ;
  SPACING 0.021 ;
  WIDTH 0.021 ;
  ENCLOSURE BELOW 0.005 0 ;
  ENCLOSURE ABOVE 0.005 0 ;
END V4

LAYER M5
  TYPE ROUTING ;
  SPACING 0.021 ;
  SPACING 0.021 SAMENET ;
  WIDTH 0.021 ;
  PITCH 0.042 ;
  AREA 0.000882 ;
  MINSIZE 0.021 0.042 ;
  DIRECTION VERTICAL ;
  PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.022 EXTENSION 0 0 0.030 ;" ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER CORNERTOCORNER WIDTH 0.000 SPACING 0.024 ; " ;
  PROPERTY LEF58_RECTONLY "RECTONLY ;" ;
END M5

LAYER V5
  TYPE CUT ;
  SPACING 0.021 ;
  WIDTH 0.021 ;
  ENCLOSURE BELOW 0.006 0 ;
  ENCLOSURE ABOVE 0.006 0 ;
END V5

LAYER M6
  TYPE ROUTING ;
  SPACING 0.038 ;
  SPACING 0.038 SAMENET ;
  WIDTH 0.038 ;
  PITCH 0.076 ;
  AREA 0.002166 ;
  MINSIZE 0.057 0.038 ;
  DIRECTION HORIZONTAL ;
  PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.039 EXTENSION 0 0 0.055 ;" ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER CORNERTOCORNER WIDTH 0.000 SPACING 0.045 ; " ;
  PROPERTY LEF58_RECTONLY "RECTONLY ;" ;
END M6

LAYER V6
  TYPE CUT ;
  SPACING 0.038 ;
  WIDTH 0.038 ;
  ENCLOSURE BELOW 0.008 0 ;
  ENCLOSURE ABOVE 0.008 0 ;
END V6

LAYER M7
  TYPE ROUTING ;
  SPACING 0.038 ;
  SPACING 0.038 SAMENET ;
  WIDTH 0.038 ;
  PITCH 0.076 ;
  AREA 0.002166 ;
  MINSIZE 0.038 0.057 ;
  DIRECTION VERTICAL ;
  PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.039 EXTENSION 0 0 0.055 ;" ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER CORNERTOCORNER WIDTH 0.000 SPACING 0.045 ; " ;
  PROPERTY LEF58_RECTONLY "RECTONLY ;" ;
END M7

LAYER V7
  TYPE CUT ;
  SPACING 0.038 ;
  WIDTH 0.038 ;
  ENCLOSURE BELOW 0.008 0 ;
  ENCLOSURE ABOVE 0.008 0 ;
END V7

LAYER M8
  TYPE ROUTING ;
  SPACING 0.038 ;
  SPACING 0.038 SAMENET ;
  WIDTH 0.038 ;
  PITCH 0.076 ;
  AREA 0.002166 ;
  MINSIZE 0.057 0.038 ;
  DIRECTION HORIZONTAL ;
  PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.039 EXTENSION 0 0 0.055 ;" ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER CORNERTOCORNER WIDTH 0.000 SPACING 0.045 ; " ;
  PROPERTY LEF58_RECTONLY "RECTONLY ;" ;
END M8

LAYER V8
  TYPE CUT ;
  SPACING 0.038 ;
  WIDTH 0.038 ;
  ENCLOSURE BELOW 0.008 0 ;
  ENCLOSURE ABOVE 0.008 0 ;
END V8

LAYER M9
  TYPE ROUTING ;
  SPACING 0.038 ;
  WIDTH 0.038 ;
  PITCH 0.076 ;
  AREA 0.002166 ;
  MINSIZE 0.038 0.057 ;
  DIRECTION VERTICAL ;
  PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.039 EXTENSION 0 0 0.055 ;" ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER CORNERTOCORNER WIDTH 0.000 SPACING 0.045 ; " ;
  PROPERTY LEF58_RECTONLY "RECTONLY ;" ;
END M9

LAYER V9
  TYPE CUT ;
  SPACING 0.038 ;
  WIDTH 0.038 ;
END V9

LAYER M10
  TYPE ROUTING ;
  SPACING 0.056 ;
  WIDTH 0.056 ;
  PITCH 0.112 ;
  DIRECTION HORIZONTAL ;
  PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.057 EXTENSION 0 0 0.080 ;" ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER CORNERTOCORNER WIDTH 0.000 SPACING 0.066 ; " ;
  PROPERTY LEF58_RECTONLY "RECTONLY ;" ;
END M10

LAYER V10
  TYPE CUT ;
  SPACING 0.056 ;
  WIDTH 0.056 ;
END V10

LAYER M11
  TYPE ROUTING ;
  SPACING 0.056 ;
  WIDTH 0.056 ;
  PITCH 0.112 ;
  DIRECTION VERTICAL ;
  PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.057 EXTENSION 0 0 0.080 ;" ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER CORNERTOCORNER WIDTH 0.000 SPACING 0.066 ; " ;
  PROPERTY LEF58_RECTONLY "RECTONLY ;" ;
END M11

LAYER V11
  TYPE CUT ;
  SPACING 0.056 ;
  WIDTH 0.056 ;
END V11

LAYER M12
  TYPE ROUTING ;
  SPACING 0.36 ;
  WIDTH 0.36 ;
  PITCH 0.72 ;
  DIRECTION HORIZONTAL ;
  PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.361 EXTENSION 0 0 0.450 ;" ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER CORNERTOCORNER WIDTH 0.000 SPACING 0.450 ; " ;
  PROPERTY LEF58_RECTONLY "RECTONLY ;" ;
END M12

LAYER V12
  TYPE CUT ;
  SPACING 0.056 ;
  WIDTH 0.056 ;
END V12

LAYER M13
  TYPE ROUTING ;
  SPACING 0.36 ;
  WIDTH 0.36 ;
  PITCH 0.72 ;
  DIRECTION VERTICAL ;
  PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.361 EXTENSION 0 0 0.450 ;" ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER CORNERTOCORNER WIDTH 0.000 SPACING 0.450 ; " ;
  PROPERTY LEF58_RECTONLY "RECTONLY ;" ;
END M13

LAYER V13
  TYPE CUT ;
  SPACING 0.056 ;
  WIDTH 0.056 ;
END V13

LAYER RDL
  TYPE ROUTING ;
  SPACING 1.6 ;
  WIDTH 1.6 ;
  PITCH 3.2 ;
  DIRECTION HORIZONTAL ;
END RDL

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP


VIA V0_0 DEFAULT
  LAYER V0 ;
    RECT -0.007 -0.006 0.007 0.006 ;
  LAYER M0 ;
    RECT -0.011 -0.006 0.011 0.006 ;
  LAYER M1 ;
    RECT -0.007 -0.010 0.007 0.010 ;
END V0_0

VIA V1_0 DEFAULT
  LAYER V1 ;
    RECT -0.007 -0.006 0.007 0.006 ;
  LAYER M1 ;
    RECT -0.007 -0.010 0.007 0.010 ;
  LAYER M2 ;
    RECT -0.011 -0.006 0.011 0.006 ;
END V1_0

VIA V2_0 DEFAULT
  LAYER V2 ;
    RECT -0.007 -0.006 0.007 0.006 ;
  LAYER M2 ;
    RECT -0.011 -0.006 0.011 0.006 ;
  LAYER M3 ;
    RECT -0.007 -0.010 0.007 0.010 ;
END V2_0

VIA V3_0 DEFAULT
  LAYER V3 ;
    RECT -0.007 -0.0105 0.007 0.0105 ;
  LAYER M3 ;
    RECT -0.007 -0.0145 0.007 0.0145 ;
  LAYER M4 ;
    RECT -0.011 -0.0105 0.011 0.0105 ;
END V3_0

VIA V4_0 DEFAULT
  LAYER V4 ;
    RECT -0.0105 -0.0105 0.0105 0.0105 ;
  LAYER M4 ;
    RECT -0.0155 -0.0105 0.0155 0.0105 ;
  LAYER M5 ;
    RECT -0.0105	-0.0155	0.0105	0.0155 ;
END V4_0

VIA V5_0 DEFAULT
  LAYER V5 ;
    RECT  -0.0105	-0.019	0.0105	0.019 ;
  LAYER M5 ;
    RECT -0.0105	-0.025	0.0105	0.025 ;
  LAYER M6 ;
    RECT -0.0165	-0.019	0.0165	0.019 ;
END V5_0

VIA V6_0 DEFAULT
  LAYER V6 ;
    RECT -0.0190	-0.0190	0.0190	0.0190 ;
  LAYER M6 ;
    RECT -0.0270	-0.0190	0.0270	0.0190 ;
  LAYER M7 ;
    RECT -0.0190	-0.0270	0.0190	0.0270 ;
END V6_0

VIA V7_0 DEFAULT
  LAYER V7 ;
    RECT -0.019	-0.019	0.019	0.019 ;
  LAYER M7 ;
    RECT -0.019	-0.027	0.019	0.027 ;
  LAYER M8 ;
    RECT -0.027	-0.019	0.027	0.019 ;
END V7_0

VIA V8_0 DEFAULT
  LAYER V8 ;
    RECT -0.0190	-0.0190	0.0190	0.0190 ;
  LAYER M8 ;
    RECT -0.0270	-0.0190	0.0270	0.0190 ;
  LAYER M9 ;
    RECT -0.0190	-0.0270	0.0190	0.0270 ;
END V8_0

VIA V9_0 DEFAULT
  LAYER V9 ;
    RECT -0.019	-0.028	0.019	0.028 ;
  LAYER M9 ;
    RECT -0.019	-0.038	0.019	0.038 ;
  LAYER M10 ;
    RECT -0.029	-0.028	0.029	0.028 ;
END V9_0

VIA V10_0 DEFAULT
  LAYER V10 ;
    RECT -0.0280	-0.0280	0.0280	0.0280 ;
  LAYER M10 ;
    RECT -0.0400	-0.0280	0.0400	0.0280 ;
  LAYER M11 ;
    RECT -0.0280	-0.0400	0.0280	0.0400 ;
END V10_0

VIA V11_0 DEFAULT
  LAYER V11 ;
    RECT -0.028	-0.18	0.028	0.18 ;
  LAYER M11 ;
    RECT -0.028	-0.192	0.028	0.192 ;
  LAYER M12 ;
    RECT -0.04	-0.18	0.04	0.18 ;
END V11_0

VIA V12_0 DEFAULT
  LAYER V12 ;
    RECT -0.1800	-0.1800	0.1800	0.1800 ;
  LAYER M12 ;
    RECT -0.2000	-0.1800	0.2000	0.1800 ;
  LAYER M13 ;
    RECT -0.1800	-0.2000	0.1800	0.2000 ;
END V12_0

VIA V13_0 DEFAULT
  LAYER V13 ;
    RECT -0.18	-0.8	0.18	0.8 ;
  LAYER M13 ;
    RECT -0.18	-0.84	0.18	0.84 ;
  LAYER RDL ;
    RECT -0.38	-0.8	0.38	0.8 ;
END V13_0

VIARULE Via0Array GENERATE
  LAYER M0 ;
    ENCLOSURE 0.004 0 ;
  LAYER M1 ;
    ENCLOSURE 0 0.004 ;
  LAYER V0 ;
    RECT -0.007 -0.006 0.007 0.006 ;
    SPACING 0.014 BY 0.012 ;
END Via0Array

VIARULE Via1Array GENERATE
  LAYER M1 ;
    ENCLOSURE 0 0.004 ;
  LAYER M2 ;
    ENCLOSURE 0.004 0 ;
  LAYER V1 ;
    RECT -0.007 -0.006 0.007 0.006 ;
    SPACING 0.028 BY 0.024 ;
END Via1Array

VIARULE Via2Array GENERATE
  LAYER M2 ;
    ENCLOSURE 0.004 0 ;
  LAYER M3 ;
    ENCLOSURE 0 0.004 ;
  LAYER V2 ;
    RECT -0.007 -0.006 0.007 0.006 ;
    SPACING 0.028 BY 0.024 ;
END Via2Array

VIARULE Via3Array GENERATE
  LAYER M3 ;
    ENCLOSURE 0 0.004 ;
  LAYER M4 ;
    ENCLOSURE 0.004 0 ;
  LAYER V3 ;
    RECT -0.007 -0.0105 0.007 0.0105 ;
    SPACING 0.028 BY 0.042 ;
END Via3Array

VIARULE Via4Array GENERATE
  LAYER M4 ;
    ENCLOSURE 0.005 0 ;
  LAYER M5 ;
    ENCLOSURE 0 0.005 ;
  LAYER V4 ;
    RECT -0.0105 -0.105 0.0105 0.0105 ;
    SPACING 0.042 BY 0.042 ;
END Via4Array

VIARULE Via5Array GENERATE
  LAYER M5 ;
    ENCLOSURE 0 0.006 ;
  LAYER M6 ;
    ENCLOSURE 0.006 0 ;
  LAYER V5 ;
    RECT -0.0105 -0.019 0.0105 0.019 ;
    SPACING 0.042 BY 0.076 ;
END Via5Array

VIARULE Via6Array GENERATE
  LAYER M6 ;
    ENCLOSURE 0.008 0 ;
  LAYER M7 ;
    ENCLOSURE 0 0.008 ;
  LAYER V6 ;
    RECT -0.019 -0.019 0.019 0.019 ;
    SPACING 0.076 BY 0.076 ;
END Via6Array

VIARULE Via7Array GENERATE
  LAYER M7 ;
    ENCLOSURE 0 0.008 ;
  LAYER M8 ;
    ENCLOSURE 0.008 0 ;
  LAYER V7 ;
    RECT -0.019 -0.019 0.019 0.019 ;
    SPACING 0.076 BY 0.076 ;
END Via7Array

VIARULE Via8Array GENERATE
  LAYER M8 ;
    ENCLOSURE 0.008 0 ;
  LAYER M9 ;
    ENCLOSURE 0 0.008 ;
  LAYER V8 ;
    RECT -0.019 -0.019 0.019 0.019  ;
    SPACING 0.076 BY 0.076 ;
END Via8Array

VIARULE Via9Array GENERATE
  LAYER M9 ;
    ENCLOSURE 0 0.010 ;
  LAYER M10 ;
    ENCLOSURE 0.010 0 ;
  LAYER V9 ;
    RECT -0.019 -0.028 0.019 0.028 ;
    SPACING 0.076 BY 0.112 ;
END Via9Array

VIARULE Via10Array GENERATE
  LAYER M10 ;
    ENCLOSURE 0.012 0 ;
  LAYER M11 ;
    ENCLOSURE 0 0.012 ;
  LAYER V10 ;
    RECT -0.028 -0.028 0.028 0.028 ;
    SPACING 0.112 BY 0.112 ;
END Via10Array

VIARULE Via11Array GENERATE
  LAYER M11 ;
    ENCLOSURE 0 0.012 ;
  LAYER M12 ;
    ENCLOSURE 0.012 0 ;
  LAYER V11 ;
    RECT -0.028 -0.18 0.028 0.18 ;
    SPACING 0.112 BY 0.72 ;
END Via11Array

VIARULE Via12Array GENERATE
  LAYER M12 ;
    ENCLOSURE 0.020 0 ;
  LAYER M13 ;
    ENCLOSURE 0 0.020 ;
  LAYER V12 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    SPACING 0.72 BY 0.72 ;
END Via12Array

VIARULE Via13Array GENERATE
  LAYER M13 ;
    ENCLOSURE 0 0.04 ;
  LAYER RDL ;
    ENCLOSURE 0.2 0 ;
  LAYER V13 ;
    RECT -0.18 -0.8 0.18 0.8 ;
    SPACING 0.72 BY 3.2 ;
END Via13Array


END LIBRARY

